///////////////////////////////////////////////////////////////////////////
// Engineer: Pietro Alberto Levo
// File: PCinc.v
// Description: implementation of the PC incrementer (adder of 4) 
///////////////////////////////////////////////////////////////////////////

module PCinc (pcOut, pcNew);
	input		[31:0] pcOut;
	output	[31:0] pcNew;
	
	assign pcNew = pcOut + 4;
	
endmodule